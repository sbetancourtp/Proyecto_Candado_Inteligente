`define B115200 868

`define B9600   10417


